module dumb_cs( //choose single chars or nums or signals
	input             clock_sink_clk,         //    clock_sink.clk
	input             reset_sink_reset,       //    reset_sink.reset
    input  [5:0]      select,
    output [15:0]     n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
);

reg [15:0] num[23:0];
assign n0 = num[0];
assign n1 = num[1];
assign n2 = num[2];
assign n3 = num[3];
assign n4 = num[4];
assign n5 = num[5];
assign n6 = num[6];
assign n7 = num[7];
assign n8 = num[8];
assign n9 = num[9];
assign n10 = num[10];
assign n11 = num[11];
assign n12 = num[12];
assign n13 = num[13];
assign n14 = num[14];
assign n15 = num[15];
assign n16 = num[16];
assign n17 = num[17];
assign n18 = num[18];
assign n19 = num[19];
assign n20 = num[20];
assign n21 = num[21];
assign n22 = num[22];
assign n23 = num[23];

always @(posedge clock_sink_clk)begin
    if(reset_sink_reset)begin
                num[0]<=16'h0000;
                num[1]<=16'h0000;
                num[2]<=16'h0000;
                num[3]<=16'h0000;
                num[4]<=16'h0000;
                num[5]<=16'h0000;
                num[6]<=16'h0000;
                num[7]<=16'h0000;
                num[8]<=16'h0000;
                num[9]<=16'h0000;
                num[10]<=16'h0000;
                num[11]<=16'h0000;
                num[12]<=16'h0000;
                num[13]<=16'h0000;
                num[14]<=16'h0000;
                num[15]<=16'h0000;
                num[16]<=16'h0000;
                num[17]<=16'h0000;
                num[18]<=16'h0000;
                num[19]<=16'h0000;
                num[20]<=16'h0000;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
    end else begin
        case (select)
            6'd0: begin
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h07E0;
                num[5] <=16'h0FF0;
                num[6] <=16'h1C38;
                num[7] <=16'h3C3C;
                num[8] <=16'h781C;
                num[9] <=16'h781E;
                num[10]<=16'h781E;
                num[11]<=16'h781E;
                num[12]<=16'h781E;
                num[13]<=16'h781E;
                num[14]<=16'h781E;
                num[15]<=16'h781E;
                num[16]<=16'h781E;
                num[17]<=16'h383C;
                num[18]<=16'h3C38;
                num[19]<=16'h1E78;
                num[20]<=16'h07E0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd1: begin
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h00C0;
                num[5] <=16'h0FC0;
                num[6] <=16'h1FC0;
                num[7] <=16'h03C0;
                num[8] <=16'h03C0;
                num[9] <=16'h03C0;
                num[10]<=16'h03C0;
                num[11]<=16'h03C0;
                num[12]<=16'h03C0;
                num[13]<=16'h03C0;
                num[14]<=16'h03C0;
                num[15]<=16'h03C0;
                num[16]<=16'h03C0;
                num[17]<=16'h03C0;
                num[18]<=16'h03C0;
                num[19]<=16'h03E0;
                num[20]<=16'h1FFC;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd2:begin
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h07E0;
                num[5] <=16'h1EF8;
                num[6] <=16'h383C;
                num[7] <=16'h781C;
                num[8] <=16'h7C1C;
                num[9] <=16'h381C;
                num[10]<=16'h003C;
                num[11]<=16'h0038;
                num[12]<=16'h0070;
                num[13]<=16'h01E0;
                num[14]<=16'h0380;
                num[15]<=16'h0700;
                num[16]<=16'h0E06;
                num[17]<=16'h1C0E;
                num[18]<=16'h301C;
                num[19]<=16'h7FFC;
                num[20]<=16'h7FFC;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end 
            6'd3:  begin
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h07E0;
                num[5] <=16'h1EF0;
                num[6] <=16'h3838;
                num[7] <=16'h383C;
                num[8] <=16'h383C;
                num[9] <=16'h003C;
                num[10]<=16'h0078;
                num[11]<=16'h03F0;
                num[12]<=16'h03F0;
                num[13]<=16'h0038;
                num[14]<=16'h001C;
                num[15]<=16'h001E;
                num[16]<=16'h381E;
                num[17]<=16'h781E;
                num[18]<=16'h783C;
                num[19]<=16'h3C78;
                num[20]<=16'h0FE0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd4: begin
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h0070;
                num[5] <=16'h0070;
                num[6] <=16'h00F0;
                num[7] <=16'h01F0;
                num[8] <=16'h03F0;
                num[9] <=16'h0770;
                num[10]<=16'h0E70;
                num[11]<=16'h0C70;
                num[12]<=16'h1870;
                num[13]<=16'h3070;
                num[14]<=16'h7070;
                num[15]<=16'hFFFF;
                num[16]<=16'h0070;
                num[17]<=16'h0070;
                num[18]<=16'h0070;
                num[19]<=16'h00F8;
                num[20]<=16'h07FE;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd5: begin
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h1FFC;
                num[5] <=16'h1FFC;
                num[6] <=16'h3800;
                num[7] <=16'h3800;
                num[8] <=16'h3800;
                num[9] <=16'h3800;
                num[10]<=16'h3FF0;
                num[11]<=16'h3FF8;
                num[12]<=16'h383C;
                num[13]<=16'h101C;
                num[14]<=16'h001E;
                num[15]<=16'h001E;
                num[16]<=16'h381E;
                num[17]<=16'h781C;
                num[18]<=16'h783C;
                num[19]<=16'h3C78;
                num[20]<=16'h0FF0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd6:begin
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h03F0;
                num[5] <=16'h0F38;
                num[6] <=16'h1C3C;
                num[7] <=16'h383C;
                num[8] <=16'h3800;
                num[9] <=16'h7800;
                num[10]<=16'h7BF0;
                num[11]<=16'h7FF8;
                num[12]<=16'h7C3C;
                num[13]<=16'h781E;
                num[14]<=16'h781E;
                num[15]<=16'h781E;
                num[16]<=16'h781E;
                num[17]<=16'h381E;
                num[18]<=16'h3C1C;
                num[19]<=16'h1E38;
                num[20]<=16'h07F0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd7: begin
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h3FFE;
                num[5] <=16'h3FFE;
                num[6] <=16'h381C;
                num[7] <=16'h7018;
                num[8] <=16'h7030;
                num[9] <=16'h0070;
                num[10]<=16'h00E0;
                num[11]<=16'h00E0;
                num[12]<=16'h01C0;
                num[13]<=16'h01C0;
                num[14]<=16'h0380;
                num[15]<=16'h0380;
                num[16]<=16'h0780;
                num[17]<=16'h0780;
                num[18]<=16'h0780;
                num[19]<=16'h0780;
                num[20]<=16'h0780;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd8: begin
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h07E0;
                num[5] <=16'h1E78;
                num[6] <=16'h381C;
                num[7] <=16'h701E;
                num[8] <=16'h701E;
                num[9] <=16'h781C;
                num[10]<=16'h3E3C;
                num[11]<=16'h1FF0;
                num[12]<=16'h1FF0;
                num[13]<=16'h3CF8;
                num[14]<=16'h783C;
                num[15]<=16'h701E;
                num[16]<=16'h701E;
                num[17]<=16'h701E;
                num[18]<=16'h701C;
                num[19]<=16'h3C38;
                num[20]<=16'h0FF0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd9: begin
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h0FE0;
                num[5] <=16'h1EF8;
                num[6] <=16'h3838;
                num[7] <=16'h781C;
                num[8] <=16'h701E;
                num[9] <=16'h701E;
                num[10]<=16'h701E;
                num[11]<=16'h781E;
                num[12]<=16'h783E;
                num[13]<=16'h3FFE;
                num[14]<=16'h0FDE;
                num[15]<=16'h001C;
                num[16]<=16'h003C;
                num[17]<=16'h1838;
                num[18]<=16'h3C78;
                num[19]<=16'h3CF0;
                num[20]<=16'h1FC0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end                     //numbers end
            6'd10: begin            //A
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h03C0;
                num[5] <=16'h03C0;
                num[6] <=16'h03C0;
                num[7] <=16'h07E0;
                num[8] <=16'h07E0;
                num[9] <=16'h0EE0;
                num[10]<=16'h0EF0;
                num[11]<=16'h0CF0;
                num[12]<=16'h1C70;
                num[13]<=16'h1C70;
                num[14]<=16'h1FF8;
                num[15]<=16'h3838;
                num[16]<=16'h3838;
                num[17]<=16'h303C;
                num[18]<=16'h701C;
                num[19]<=16'h701E;
                num[20]<=16'hFC7F;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd11: begin            //B
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'hFFE0;
                num[5] <=16'h7FF8;
                num[6] <=16'h383C;
                num[7] <=16'h381E;
                num[8] <=16'h381E;
                num[9] <=16'h381C;
                num[10]<=16'h383C;
                num[11]<=16'h3FF8;
                num[12]<=16'h3FF8;
                num[13]<=16'h381C;
                num[14]<=16'h381E;
                num[15]<=16'h380F;
                num[16]<=16'h380F;
                num[17]<=16'h380E;
                num[18]<=16'h381E;
                num[19]<=16'h387C;
                num[20]<=16'hFFF0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd12: begin            //C
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h03FE;
                num[5] <=16'h0F3E;
                num[6] <=16'h1C0E;
                num[7] <=16'h3806;
                num[8] <=16'h7807;
                num[9] <=16'h7800;
                num[10]<=16'hF000;
                num[11]<=16'hF000;
                num[12]<=16'hF000;
                num[13]<=16'hF000;
                num[14]<=16'hF000;
                num[15]<=16'h7000;
                num[16]<=16'h7807;
                num[17]<=16'h7806;
                num[18]<=16'h3C0C;
                num[19]<=16'h1F3C;
                num[20]<=16'h07F0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd13: begin            //D
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'hFF80;
                num[5] <=16'h7FF0;
                num[6] <=16'h3838;
                num[7] <=16'h381C;
                num[8] <=16'h381E;
                num[9] <=16'h381E;
                num[10]<=16'h380E;
                num[11]<=16'h380F;
                num[12]<=16'h380F;
                num[13]<=16'h380F;
                num[14]<=16'h380E;
                num[15]<=16'h381E;
                num[16]<=16'h381E;
                num[17]<=16'h381C;
                num[18]<=16'h383C;
                num[19]<=16'h38F0;
                num[20]<=16'hFFC0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd14: begin            //E
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'hFFFC;
                num[5] <=16'h7FFC;
                num[6] <=16'h3C0E;
                num[7] <=16'h3C06;
                num[8] <=16'h3C00;
                num[9] <=16'h3C30;
                num[10]<=16'h3C30;
                num[11]<=16'h3FF0;
                num[12]<=16'h3FF0;
                num[13]<=16'h3C30;
                num[14]<=16'h3C30;
                num[15]<=16'h3C00;
                num[16]<=16'h3C00;
                num[17]<=16'h3C07;
                num[18]<=16'h3C0E;
                num[19]<=16'h3C1E;
                num[20]<=16'hFFFC;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd15: begin            //F
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'hFFFE;
                num[5] <=16'h7FFE;
                num[6] <=16'h3C0E;
                num[7] <=16'h3C07;
                num[8] <=16'h3C00;
                num[9] <=16'h3C18;
                num[10]<=16'h3C38;
                num[11]<=16'h3C78;
                num[12]<=16'h3FF8;
                num[13]<=16'h3C38;
                num[14]<=16'h3C38;
                num[15]<=16'h3C00;
                num[16]<=16'h3C00;
                num[17]<=16'h3C00;
                num[18]<=16'h3C00;
                num[19]<=16'h3C00;
                num[20]<=16'hFF00;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd16: begin            //G
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h07F8;
                num[5] <=16'h0F7C;
                num[6] <=16'h1C1C;
                num[7] <=16'h381C;
                num[8] <=16'h780C;
                num[9] <=16'h7000;
                num[10]<=16'hF000;
                num[11]<=16'hF000;
                num[12]<=16'hF000;
                num[13]<=16'hF07F;
                num[14]<=16'hF07E;
                num[15]<=16'hF01C;
                num[16]<=16'h701C;
                num[17]<=16'h781C;
                num[18]<=16'h381C;
                num[19]<=16'h1E3C;
                num[20]<=16'h0FF0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd17: begin            //H
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'hFC7F;
                num[5] <=16'h7C3E;
                num[6] <=16'h781C;
                num[7] <=16'h781C;
                num[8] <=16'h781C;
                num[9] <=16'h781C;
                num[10]<=16'h781C;
                num[11]<=16'h781C;
                num[12]<=16'h7FFC;
                num[13]<=16'h781C;
                num[14]<=16'h781C;
                num[15]<=16'h781C;
                num[16]<=16'h781C;
                num[17]<=16'h781C;
                num[18]<=16'h781C;
                num[19]<=16'h781C;
                num[20]<=16'hFE7F;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd18: begin            //I
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h3FFC;
                num[5] <=16'h1FF8;
                num[6] <=16'h03C0;
                num[7] <=16'h03C0;
                num[8] <=16'h03C0;
                num[9] <=16'h03C0;
                num[10]<=16'h03C0;
                num[11]<=16'h03C0;
                num[12]<=16'h03C0;
                num[13]<=16'h03C0;
                num[14]<=16'h03C0;
                num[15]<=16'h03C0;
                num[16]<=16'h03C0;
                num[17]<=16'h03C0;
                num[18]<=16'h03C0;
                num[19]<=16'h03C0;
                num[20]<=16'h3FFC;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd19: begin            //J
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h0FFF;
                num[5] <=16'h07FE;
                num[6] <=16'h00F0;
                num[7] <=16'h00F0;
                num[8] <=16'h00F0;
                num[9] <=16'h00F0;
                num[10]<=16'h00F0;
                num[11]<=16'h00F0;
                num[12]<=16'h00F0;
                num[13]<=16'h00F0;
                num[14]<=16'h00F0;
                num[15]<=16'h00F0;
                num[16]<=16'h00F0;
                num[17]<=16'h00F0;
                num[18]<=16'h00F0;
                num[19]<=16'h00F0;
                num[20]<=16'h70F0;
                num[21]<=16'hF8E0;
                num[22]<=16'h7BC0;
                num[23]<=16'h3F00;
            end
            6'd20: begin            //K
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'hFE7E;
                num[5] <=16'h7E7E;
                num[6] <=16'h3838;
                num[7] <=16'h3860;
                num[8] <=16'h38E0;
                num[9] <=16'h39C0;
                num[10]<=16'h3B80;
                num[11]<=16'h3F80;
                num[12]<=16'h3FC0;
                num[13]<=16'h3DE0;
                num[14]<=16'h38E0;
                num[15]<=16'h38F0;
                num[16]<=16'h3870;
                num[17]<=16'h3878;
                num[18]<=16'h383C;
                num[19]<=16'h383E;
                num[20]<=16'hFE7F;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd21: begin            //L
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h7F00;
                num[5] <=16'h7E00;
                num[6] <=16'h3C00;
                num[7] <=16'h3C00;
                num[8] <=16'h3C00;
                num[9] <=16'h3C00;
                num[10]<=16'h3C00;
                num[11]<=16'h3C00;
                num[12]<=16'h3C00;
                num[13]<=16'h3C00;
                num[14]<=16'h3C00;
                num[15]<=16'h3C00;
                num[16]<=16'h3C00;
                num[17]<=16'h3C07;
                num[18]<=16'h3C06;
                num[19]<=16'h3C1E;
                num[20]<=16'hFFFE;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd22: begin            //M
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'hF01F;
                num[5] <=16'hF81F;
                num[6] <=16'h783E;
                num[7] <=16'h783E;
                num[8] <=16'h7C3E;
                num[9] <=16'h7C7E;
                num[10]<=16'h7C7E;
                num[11]<=16'h7E7E;
                num[12]<=16'h6EFE;
                num[13]<=16'h6EDE;
                num[14]<=16'h6EDE;
                num[15]<=16'h67DE;
                num[16]<=16'h67DE;
                num[17]<=16'h679E;
                num[18]<=16'h679E;
                num[19]<=16'h639E;
                num[20]<=16'hFB7F;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd23: begin            //N
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'hF83F;
                num[5] <=16'hFC1F;
                num[6] <=16'h3C0C;
                num[7] <=16'h3E0C;
                num[8] <=16'h3F0C;
                num[9] <=16'h370C;
                num[10]<=16'h378C;
                num[11]<=16'h33CC;
                num[12]<=16'h31CC;
                num[13]<=16'h31EC;
                num[14]<=16'h30FC;
                num[15]<=16'h307C;
                num[16]<=16'h307C;
                num[17]<=16'h303C;
                num[18]<=16'h301C;
                num[19]<=16'h301C;
                num[20]<=16'hFC0C;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd24: begin            //O
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h07E0;
                num[5] <=16'h1F78;
                num[6] <=16'h3C1C;
                num[7] <=16'h381C;
                num[8] <=16'h781E;
                num[9] <=16'h780E;
                num[10]<=16'h700F;
                num[11]<=16'hF00F;
                num[12]<=16'hF00F;
                num[13]<=16'hF00F;
                num[14]<=16'h700F;
                num[15]<=16'h700F;
                num[16]<=16'h780E;
                num[17]<=16'h381E;
                num[18]<=16'h3C1C;
                num[19]<=16'h1E78;
                num[20]<=16'h07F0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd25: begin            //P
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'hFFE0;
                num[5] <=16'h7FFC;
                num[6] <=16'h3C1E;
                num[7] <=16'h3C0E;
                num[8] <=16'h3C0E;
                num[9] <=16'h3C0E;
                num[10]<=16'h3C0E;
                num[11]<=16'h3C3C;
                num[12]<=16'h3FF8;
                num[13]<=16'h3F80;
                num[14]<=16'h3C00;
                num[15]<=16'h3C00;
                num[16]<=16'h3C00;
                num[17]<=16'h3C00;
                num[18]<=16'h3C00;
                num[19]<=16'h3C00;
                num[20]<=16'hFF00;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd26: begin            //Q
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h07E0;
                num[5] <=16'h1E78;
                num[6] <=16'h3C3C;
                num[7] <=16'h781E;
                num[8] <=16'h781E;
                num[9] <=16'h700E;
                num[10]<=16'hF00F;
                num[11]<=16'hF00F;
                num[12]<=16'hF00F;
                num[13]<=16'hF00F;
                num[14]<=16'hF00F;
                num[15]<=16'h730E;
                num[16]<=16'h7FCE;
                num[17]<=16'h7DFE;
                num[18]<=16'h3CFC;
                num[19]<=16'h1EF8;
                num[20]<=16'h07F6;
                num[21]<=16'h007E;
                num[22]<=16'h003C;
                num[23]<=16'h0000;
            end
            6'd27: begin            //R
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'hFFE0;
                num[5] <=16'h7FF8;
                num[6] <=16'h3C1C;
                num[7] <=16'h3C1E;
                num[8] <=16'h3C1E;
                num[9] <=16'h3C1E;
                num[10]<=16'h3C1C;
                num[11]<=16'h3C78;
                num[12]<=16'h3FE0;
                num[13]<=16'h3DE0;
                num[14]<=16'h3CE0;
                num[15]<=16'h3C70;
                num[16]<=16'h3C78;
                num[17]<=16'h3C38;
                num[18]<=16'h3C3C;
                num[19]<=16'h3C1C;
                num[20]<=16'hFF1F;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd28: begin            //S
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h0FE8;
                num[5] <=16'h1EFC;
                num[6] <=16'h383C;
                num[7] <=16'h701C;
                num[8] <=16'h700C;
                num[9] <=16'h7800;
                num[10]<=16'h3E00;
                num[11]<=16'h1F80;
                num[12]<=16'h07F0;
                num[13]<=16'h00F8;
                num[14]<=16'h003C;
                num[15]<=16'h001E;
                num[16]<=16'h600E;
                num[17]<=16'h700E;
                num[18]<=16'h701C;
                num[19]<=16'h7C38;
                num[20]<=16'h3FF0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000; 
            end
            6'd29: begin            //T
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h7FFC;
                num[5] <=16'h7FFE;
                num[6] <=16'h63C6;
                num[7] <=16'hE3C6;
                num[8] <=16'h43C0;
                num[9] <=16'h03C0;
                num[10]<=16'h03C0;
                num[11]<=16'h03C0;
                num[12]<=16'h03C0;
                num[13]<=16'h03C0;
                num[14]<=16'h03C0;
                num[15]<=16'h03C0;
                num[16]<=16'h03C0;
                num[17]<=16'h03C0;
                num[18]<=16'h03C0;
                num[19]<=16'h03C0;
                num[20]<=16'h0FF0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd30: begin            //U
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'hFE3F;
                num[5] <=16'hFC1E;
                num[6] <=16'h780C;
                num[7] <=16'h780C;
                num[8] <=16'h780C;
                num[9] <=16'h780C;
                num[10]<=16'h780C;
                num[11]<=16'h780C;
                num[12]<=16'h780C;
                num[13]<=16'h780C;
                num[14]<=16'h780C;
                num[15]<=16'h780C;
                num[16]<=16'h780C;
                num[17]<=16'h380C;
                num[18]<=16'h381C;
                num[19]<=16'h1E78;
                num[20]<=16'h0FE0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd31: begin            //V
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'hFC3F;
                num[5] <=16'hFC1E;
                num[6] <=16'h381C;
                num[7] <=16'h3C18;
                num[8] <=16'h3C18;
                num[9] <=16'h1C38;
                num[10]<=16'h1E30;
                num[11]<=16'h1E70;
                num[12]<=16'h0E70;
                num[13]<=16'h0F60;
                num[14]<=16'h0FE0;
                num[15]<=16'h07C0;
                num[16]<=16'h07C0;
                num[17]<=16'h07C0;
                num[18]<=16'h0380;
                num[19]<=16'h0380;
                num[20]<=16'h0380;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd32: begin            //W
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'hFFFF;
                num[5] <=16'hFBCF;
                num[6] <=16'h71C6;
                num[7] <=16'h71CE;
                num[8] <=16'h79CC;
                num[9] <=16'h79CC;
                num[10]<=16'h3BEC;
                num[11]<=16'h3BFC;
                num[12]<=16'h3BFC;
                num[13]<=16'h3FF8;
                num[14]<=16'h1FF8;
                num[15]<=16'h1EF8;
                num[16]<=16'h1E78;
                num[17]<=16'h1E70;
                num[18]<=16'h1E70;
                num[19]<=16'h0C70;
                num[20]<=16'h0C70;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;   
            end
            6'd33: begin            //X
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h7E7E;
                num[5] <=16'h7C3E;
                num[6] <=16'h1C38;
                num[7] <=16'h1E30;
                num[8] <=16'h0E70;
                num[9] <=16'h0760;
                num[10]<=16'h07C0;
                num[11]<=16'h03C0;
                num[12]<=16'h03C0;
                num[13]<=16'h03C0;
                num[14]<=16'h07E0;
                num[15]<=16'h06F0;
                num[16]<=16'h0E70;
                num[17]<=16'h0C78;
                num[18]<=16'h183C;
                num[19]<=16'h383C;
                num[20]<=16'hFC7F;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd34: begin            //Y
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'hFE3F;
                num[5] <=16'h7C3E;
                num[6] <=16'h3C18;
                num[7] <=16'h1C18;
                num[8] <=16'h1E30;
                num[9] <=16'h0E30;
                num[10]<=16'h0F60;
                num[11]<=16'h07E0;
                num[12]<=16'h07C0;
                num[13]<=16'h03C0;
                num[14]<=16'h03C0;
                num[15]<=16'h03C0;
                num[16]<=16'h03C0;
                num[17]<=16'h03C0;
                num[18]<=16'h03C0;
                num[19]<=16'h03C0;
                num[20]<=16'h0FF0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd35: begin            //Z
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h1FFE;
                num[5] <=16'h3FFE;
                num[6] <=16'h383C;
                num[7] <=16'h7038;
                num[8] <=16'h0078;
                num[9] <=16'h00F0;
                num[10]<=16'h00E0;
                num[11]<=16'h01C0;
                num[12]<=16'h03C0;
                num[13]<=16'h0780;
                num[14]<=16'h0700;
                num[15]<=16'h0F00;
                num[16]<=16'h1E00;
                num[17]<=16'h1C06;
                num[18]<=16'h380E;
                num[19]<=16'h783C;
                num[20]<=16'h7FFC;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd36: begin            //.
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h0000;
                num[5] <=16'h0000;
                num[6] <=16'h0000;
                num[7] <=16'h0000;
                num[8] <=16'h0000;
                num[9] <=16'h0000;
                num[10]<=16'h0000;
                num[11]<=16'h0000;
                num[12]<=16'h0000;
                num[13]<=16'h0000;
                num[14]<=16'h0000;
                num[15]<=16'h0000;
                num[16]<=16'h0000;
                num[17]<=16'h0000;
                num[18]<=16'h3C00;
                num[19]<=16'h7E00;
                num[20]<=16'h3C00;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd37: begin            //:
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h0000;
                num[5] <=16'h0000;
                num[6] <=16'h0000;
                num[7] <=16'h0000;
                num[8] <=16'h0000;
                num[9] <=16'h0380;
                num[10]<=16'h07C0;
                num[11]<=16'h03C0;
                num[12]<=16'h0000;
                num[13]<=16'h0000;
                num[14]<=16'h0000;
                num[15]<=16'h0000;
                num[16]<=16'h0000;
                num[17]<=16'h0000;
                num[18]<=16'h03C0;
                num[19]<=16'h07C0;
                num[20]<=16'h03C0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            6'd38: begin            //!
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h03C0;
                num[5] <=16'h03C0;
                num[6] <=16'h03C0;
                num[7] <=16'h03C0;
                num[8] <=16'h03C0;
                num[9] <=16'h03C0;
                num[10]<=16'h0380;
                num[11]<=16'h0380;
                num[12]<=16'h0180;
                num[13]<=16'h0180;
                num[14]<=16'h0180;
                num[15]<=16'h0180;
                num[16]<=16'h0000;
                num[17]<=16'h0000;
                num[18]<=16'h03C0;
                num[19]<=16'h07C0;
                num[20]<=16'h03C0;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
            default: begin
                num[0] <=16'h0000;
                num[1] <=16'h0000;
                num[2] <=16'h0000;
                num[3] <=16'h0000;
                num[4] <=16'h0000;
                num[5] <=16'h0000;
                num[6] <=16'h0000;
                num[7] <=16'h0000;
                num[8] <=16'h0000;
                num[9] <=16'h0000;
                num[10]<=16'h0000;
                num[11]<=16'h0000;
                num[12]<=16'h0000;
                num[13]<=16'h0000;
                num[14]<=16'h0000;
                num[15]<=16'h0000;
                num[16]<=16'h0000;
                num[17]<=16'h0000;
                num[18]<=16'h0000;
                num[19]<=16'h0000;
                num[20]<=16'h0000;
                num[21]<=16'h0000;
                num[22]<=16'h0000;
                num[23]<=16'h0000;
            end
        endcase
    end
end


endmodule
